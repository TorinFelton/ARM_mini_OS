//Verilog HDL for "COMP22712", "CONST_clock_divide_val" "functional"


module CONST_clock_divide_val (output[15:0] value );
	assign value = 5000;

endmodule
